library verilog;
use verilog.vl_types.all;
entity TB_ii is
end TB_ii;
