library verilog;
use verilog.vl_types.all;
entity TB_oi is
end TB_oi;
